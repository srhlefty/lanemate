----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:38:39 02/18/2019 
-- Design Name: 
-- Module Name:    generate_sd_de - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity generate_sd_de is
    Port ( PCLK : in  STD_LOGIC;
           FIELD : in  STD_LOGIC;
			  HSIN : in std_logic;
           HS : out  STD_LOGIC;
			  VS : out std_logic;
           DE : out  STD_LOGIC);
end generate_sd_de;

architecture Behavioral of generate_sd_de is

	signal oldH : std_logic := '1';
	signal oldF : std_logic := '0';
	
	signal hs_out : std_logic := '1';
	signal hcount : natural range 0 to 65535 := 0;
	
	signal vs_out : std_logic := '1';
	signal vcount : natural range 0 to 65535 := 0;
	
	signal line : natural range 0 to 511 := 0;
	
	signal de_all : std_logic := '0';
	signal de_ok : std_logic := '0';
begin

	-- If I ask the 7180 for VSYNC, it gives me a tiny pulse instead of the
	-- width specified by the standard. Here I make a new pulse.
	process(PCLK) is
	begin
	if(rising_edge(PCLK)) then
		oldF <= FIELD;
		if((oldF xor FIELD) = '1') then
			vs_out <= '0';
			vcount <= 3*1716;
		else
			if(vcount = 0) then
				vs_out <= '1';
			else
				vcount <= vcount - 1;
			end if;
		end if;
	end if;
	end process;
	
	VS <= vs_out;



	-- The HSYNC generated by the 7180 is one clock, so here I stretch it
	-- to the size specified by the standard
	process(PCLK) is
	begin
	if(rising_edge(PCLK)) then
		oldH <= HSIN;
		if(HSIN = '0' and oldH = '1') then
			hs_out <= '0';
			hcount <= 1;
		else
			hcount <= hcount + 1;
			if(hcount = 124) then
				hs_out <= '1';
			end if;
		end if;

		-- track what line I'm on for DE suppression
		if((oldF xor FIELD) = '1') then
			if(FIELD = '0') then
				-- first field?
				line <= 4;
			else
				line <= 266;
			end if;
		else
			if(HSIN = '0' and oldH = '1') then
				line <= line + 1;
			end if;
		end if;
		
	end if;
	end process;
	
	HS <= hs_out;
	
	
	-- Wrap a DE around the line
	process(PCLK) is
	begin
	if(rising_edge(PCLK)) then
		if(hcount > (124+114-1) and hcount < (124+114+1440)) then
			de_all <= '1';
		else
			de_all <= '0';
		end if;
		
		if((line >= 22 and line <= 261) or (line >= 285 and line <= 524)) then
			de_ok <= '1';
		else
			de_ok <= '0';
		end if;
	end if;
	end process;
	
	DE <= de_all and de_ok;

end Behavioral;

