--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:23:02 02/19/2019
-- Design Name:   
-- Module Name:   C:/Users/Steven/Documents/Code/lanemate/firmware/src/bt656_decode_tb.vhd
-- Project Name:  firmware
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: bt656_decode
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY bt656_decode_tb IS
END bt656_decode_tb;
 
ARCHITECTURE behavior OF bt656_decode_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT bt656_decode
    PORT(
         D : IN  std_logic_vector(7 downto 0);
         CLK : IN  std_logic;
         VS : OUT  std_logic;
         HS : OUT  std_logic;
         DE : OUT  std_logic;
         DOUT : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal D : std_logic_vector(7 downto 0) := (others => '0');
   signal CLK : std_logic := '0';

 	--Outputs
   signal VS : std_logic;
   signal HS : std_logic;
   signal DE : std_logic;
   signal DOUT : std_logic_vector(7 downto 0);

	type mem_t is array(0 to 1715) of std_logic_vector(7 downto 0);
 
	signal rom : mem_t := (
		x"FF", x"00", x"00", "10010000", -- eav
x"80", x"10", x"80", x"10", -- 268 clocks alternating 80,10
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
x"80", x"10", x"80", x"10",
		x"FF", x"00", x"00", "10000000", -- sav
x"01", x"02", x"03", x"04", -- 1440 clocks of data
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04",
x"01", x"02", x"03", x"04"		
	);

	signal count : natural := 0;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: bt656_decode PORT MAP (
          D => D,
          CLK => CLK,
          VS => VS,
          HS => HS,
          DE => DE,
          DOUT => DOUT
        );

	CLK <= not CLK after 5 ns;
	
	process(CLK) is
	begin
	if(rising_edge(CLK)) then
		if(count = rom'high) then
			count <= 0;
		else
			count <= count + 1;
		end if;
		D <= rom(count);
		
	end if;
	end process;
END;
